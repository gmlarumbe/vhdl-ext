library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity block0 is
    generic (Generic0 : integer := 0;
             Generic1 : integer := 0;
             Generic2 : integer := 0);
    port (Port0 : in std_logic;
          Port1 : in std_logic;
          Port2 : in std_logic);
end entity block0;

architecture RTL of block0 is

begin  -- architecture RTL



end architecture RTL;
